** Profile: "SCHEMATIC1-hand_pdn_v2"  [ G:\My Drive\Graduate\Project\Haptic Assistance Navigation Device\PCB Design\Simulation\paper\hand_pdn_v2-pspicefiles\schematic1\hand_pdn_v2.sim ] 

** Creating circuit file "hand_pdn_v2.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../third_party/ti/tps63805/tps63805_trans.lib" 
.LIB "../../../third_party/ti/tps63806/tps63806_trans.lib" 
.LIB "../../../third_party/ti/tps61023/library/tps61023_trans.lib" 
.LIB "../../../third_party/diode inc/dmp2035uvt.lib" 
.LIB "../../../third_party/ti/tps22965/tps22965_trans.lib" 
.LIB "../../../third_party/murata/ferrite bead/blm18sg700tz1.lib" 
* From [PSPICE NETLIST] section of D:\Dennis\Develop\Simulation\ORCAD\Project\cdssetup\OrCAD_PSpice\22.1.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 35m 0.1m 2n 
.OPTIONS ADVCONV
.OPTIONS ABSTOL= 1e-9
.OPTIONS RELTOL= 0.005
.OPTIONS VNTOL= 1e-6
.OPTIONS SPEED_LEVEL= 0
.AUTOCONVERGE ITL1=1000 ITL2=1000 ITL4=1000 RELTOL=0.05 ABSTOL=1.0E-6 VNTOL=.001 PIVTOL=1.0E-10 
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
