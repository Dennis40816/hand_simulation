** Profile: "STARTUP-tran"  [ C:\Dennis\Develop\Simulation\ORCAD\Project\hand_pdn_v2\third_party\TI\TPS63806\tps63806_trans-pspicefiles\startup\tran.sim ] 

** Creating circuit file "tran.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../tps63806_trans.lib" 
* From [PSPICE NETLIST] section of C:\Dennis\Develop\Simulation\ORCAD\cdssetup\OrCAD_PSpice\22.1.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 0.45m 0 10n 
.OPTIONS ADVCONV
.OPTIONS ABSTOL= 1.0n
.OPTIONS ITL4= 30
.PROBE64 V(alias(*)) I(alias(*)) 
.INC "..\STARTUP.net" 


.END
